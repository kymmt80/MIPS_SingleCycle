module inst_mem(input [31:0]Address,output reg [31:0]inst);
reg [31:0] mem[0:1023];

initial begin
    mem[0]=32'b00100000000000010000000000101000;//addi R1 R0 36
    mem[1]=32'b00100000000001010000000000000000;//addi R5 R0 0
    mem[2]=32'b00010000001000000000000000000100;//beq R1 R0 END //LOOP
    mem[3]=32'b10001100001001000000001111100100;//lw  R4 1000(R1)
    mem[4]=32'b00000000101001000010100000100000;//add R5 R4 R5
    mem[5]=32'b00100000001000011111111111111100;//addi R1 R1 -4
    mem[6]=32'b00001000000000000000000000000010;//J LOOP
    mem[7]=32'b10101100000001010000011111010000;//sw R5 2000(R0) //END
end

always @(Address) begin
    inst<=mem[Address[31:2]];
end
endmodule